module Clock(
	input logic clock,
	output logic clock_dec,
	output logic clock_sec
); 


endmodule
